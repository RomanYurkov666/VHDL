// rangefinder_sopc.v

// Generated using ACDS version 14.0 200 at 2017.05.29.21:21:27

`timescale 1 ps / 1 ps
module rangefinder_sopc (
		input  wire       clk_clk,                           //                 clk.clk
		input  wire       reset_reset_n,                     //               reset.reset_n
		output wire       sys_timer_export,                  //           sys_timer.export
		input  wire       pc_uart_rxd,                       //             pc_uart.rxd
		output wire       pc_uart_txd,                       //                    .txd
		output wire [7:0] leds_port_export,                  //           leds_port.export
		inout  wire [1:0] i2c_port_export,                   //            i2c_port.export
		input  wire       laser_driver_ref_clk,              //        laser_driver.ref_clk
		input  wire       laser_driver_driver_enable,        //                    .driver_enable
		output wire       laser_driver_laser,                //                    .laser
		input  wire       laser_driver_comparator,           //                    .comparator
		output wire       spi_tdc_master_clk,                //             spi_tdc.master_clk
		output wire       spi_tdc_master_csn,                //                    .master_csn
		output wire       spi_tdc_master_mosi,               //                    .master_mosi
		input  wire       spi_tdc_master_miso,               //                    .master_miso
		output wire       pulse_generator_start_pulse,       //     pulse_generator.start_pulse
		output wire       pulse_generator_stop_pulse,        //                    .stop_pulse
		output wire       spi_vga_master_clk,                //             spi_vga.master_clk
		output wire       spi_vga_master_csn,                //                    .master_csn
		output wire       spi_vga_master_mosi,               //                    .master_mosi
		input  wire       spi_vga_master_miso,               //                    .master_miso
		output wire       rs485_de_export,                   //            rs485_de.export
		output wire       tdc_enable_export,                 //          tdc_enable.export
		output wire       system_mode_export,                //         system_mode.export
		output wire       amp_gain_export,                   //            amp_gain.export
		input  wire       apd_overcurrent_export,            //     apd_overcurrent.export
		output wire       spi_apd_master_clk,                //             spi_apd.master_clk
		output wire       spi_apd_master_csn,                //                    .master_csn
		output wire       spi_apd_master_mosi,               //                    .master_mosi
		input  wire       spi_apd_master_miso,               //                    .master_miso
		output wire       iris_motor_dir,                    //                iris.motor_dir
		output wire       iris_motor_step,                   //                    .motor_step
		output wire       iris_motor_en,                     //                    .motor_en
		output wire       atten_motor_dir,                   //               atten.motor_dir
		output wire       atten_motor_step,                  //                    .motor_step
		output wire       atten_motor_en,                    //                    .motor_en
		input  wire       laser_charge_ref_clk,              //        laser_charge.ref_clk
		input  wire       laser_charge_driver_enable,        //                    .driver_enable
		output wire       laser_charge_laser,                //                    .laser
		input  wire       laser_charge_comparator,           //                    .comparator
		input  wire       tdc_start_pulse_gen_ref_clk,       // tdc_start_pulse_gen.ref_clk
		input  wire       tdc_start_pulse_gen_driver_enable, //                    .driver_enable
		output wire       tdc_start_pulse_gen_laser,         //                    .laser
		input  wire       tdc_start_pulse_gen_comparator,    //                    .comparator
		input  wire       adc_clk_clk,                       //             adc_clk.clk
		input  wire [7:0] adc_data_adc_data,                 //            adc_data.adc_data
		input  wire       adc_data_comparator                //                    .comparator
	);

	wire         cpu_instruction_master_waitrequest;                              // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [15:0] cpu_instruction_master_address;                                  // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                     // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                 // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_readdatavalid;                            // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         cpu_data_master_waitrequest;                                     // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                       // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [15:0] cpu_data_master_address;                                         // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                           // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                            // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                        // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                     // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire         cpu_data_master_readdatavalid;                                   // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire   [3:0] cpu_data_master_byteenable;                                      // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;             // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;               // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                 // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                   // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                    // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;             // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;              // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_ram_cpu_s1_writedata;                          // mm_interconnect_0:ram_cpu_s1_writedata -> ram_cpu:writedata
	wire  [12:0] mm_interconnect_0_ram_cpu_s1_address;                            // mm_interconnect_0:ram_cpu_s1_address -> ram_cpu:address
	wire         mm_interconnect_0_ram_cpu_s1_chipselect;                         // mm_interconnect_0:ram_cpu_s1_chipselect -> ram_cpu:chipselect
	wire         mm_interconnect_0_ram_cpu_s1_clken;                              // mm_interconnect_0:ram_cpu_s1_clken -> ram_cpu:clken
	wire         mm_interconnect_0_ram_cpu_s1_write;                              // mm_interconnect_0:ram_cpu_s1_write -> ram_cpu:write
	wire  [31:0] mm_interconnect_0_ram_cpu_s1_readdata;                           // ram_cpu:readdata -> mm_interconnect_0:ram_cpu_s1_readdata
	wire   [3:0] mm_interconnect_0_ram_cpu_s1_byteenable;                         // mm_interconnect_0:ram_cpu_s1_byteenable -> ram_cpu:byteenable
	wire  [31:0] mm_interconnect_0_ram_cpu_s2_writedata;                          // mm_interconnect_0:ram_cpu_s2_writedata -> ram_cpu:writedata2
	wire  [12:0] mm_interconnect_0_ram_cpu_s2_address;                            // mm_interconnect_0:ram_cpu_s2_address -> ram_cpu:address2
	wire         mm_interconnect_0_ram_cpu_s2_chipselect;                         // mm_interconnect_0:ram_cpu_s2_chipselect -> ram_cpu:chipselect2
	wire         mm_interconnect_0_ram_cpu_s2_clken;                              // mm_interconnect_0:ram_cpu_s2_clken -> ram_cpu:clken2
	wire         mm_interconnect_0_ram_cpu_s2_write;                              // mm_interconnect_0:ram_cpu_s2_write -> ram_cpu:write2
	wire  [31:0] mm_interconnect_0_ram_cpu_s2_readdata;                           // ram_cpu:readdata2 -> mm_interconnect_0:ram_cpu_s2_readdata
	wire   [3:0] mm_interconnect_0_ram_cpu_s2_byteenable;                         // mm_interconnect_0:ram_cpu_s2_byteenable -> ram_cpu:byteenable2
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;                  // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;                 // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire  [15:0] mm_interconnect_0_sys_timer_s1_writedata;                        // mm_interconnect_0:sys_timer_s1_writedata -> sys_timer:writedata
	wire   [2:0] mm_interconnect_0_sys_timer_s1_address;                          // mm_interconnect_0:sys_timer_s1_address -> sys_timer:address
	wire         mm_interconnect_0_sys_timer_s1_chipselect;                       // mm_interconnect_0:sys_timer_s1_chipselect -> sys_timer:chipselect
	wire         mm_interconnect_0_sys_timer_s1_write;                            // mm_interconnect_0:sys_timer_s1_write -> sys_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_timer_s1_readdata;                         // sys_timer:readdata -> mm_interconnect_0:sys_timer_s1_readdata
	wire  [15:0] mm_interconnect_0_pc_uart_s1_writedata;                          // mm_interconnect_0:pc_uart_s1_writedata -> pc_uart:writedata
	wire   [2:0] mm_interconnect_0_pc_uart_s1_address;                            // mm_interconnect_0:pc_uart_s1_address -> pc_uart:address
	wire         mm_interconnect_0_pc_uart_s1_chipselect;                         // mm_interconnect_0:pc_uart_s1_chipselect -> pc_uart:chipselect
	wire         mm_interconnect_0_pc_uart_s1_write;                              // mm_interconnect_0:pc_uart_s1_write -> pc_uart:write_n
	wire         mm_interconnect_0_pc_uart_s1_read;                               // mm_interconnect_0:pc_uart_s1_read -> pc_uart:read_n
	wire  [15:0] mm_interconnect_0_pc_uart_s1_readdata;                           // pc_uart:readdata -> mm_interconnect_0:pc_uart_s1_readdata
	wire         mm_interconnect_0_pc_uart_s1_begintransfer;                      // mm_interconnect_0:pc_uart_s1_begintransfer -> pc_uart:begintransfer
	wire  [31:0] mm_interconnect_0_leds_port_s1_writedata;                        // mm_interconnect_0:leds_port_s1_writedata -> leds_port:writedata
	wire   [2:0] mm_interconnect_0_leds_port_s1_address;                          // mm_interconnect_0:leds_port_s1_address -> leds_port:address
	wire         mm_interconnect_0_leds_port_s1_chipselect;                       // mm_interconnect_0:leds_port_s1_chipselect -> leds_port:chipselect
	wire         mm_interconnect_0_leds_port_s1_write;                            // mm_interconnect_0:leds_port_s1_write -> leds_port:write_n
	wire  [31:0] mm_interconnect_0_leds_port_s1_readdata;                         // leds_port:readdata -> mm_interconnect_0:leds_port_s1_readdata
	wire  [31:0] mm_interconnect_0_i2c_port_s1_writedata;                         // mm_interconnect_0:i2c_port_s1_writedata -> i2c_port:writedata
	wire   [2:0] mm_interconnect_0_i2c_port_s1_address;                           // mm_interconnect_0:i2c_port_s1_address -> i2c_port:address
	wire         mm_interconnect_0_i2c_port_s1_chipselect;                        // mm_interconnect_0:i2c_port_s1_chipselect -> i2c_port:chipselect
	wire         mm_interconnect_0_i2c_port_s1_write;                             // mm_interconnect_0:i2c_port_s1_write -> i2c_port:write_n
	wire  [31:0] mm_interconnect_0_i2c_port_s1_readdata;                          // i2c_port:readdata -> mm_interconnect_0:i2c_port_s1_readdata
	wire  [31:0] mm_interconnect_0_laser_driver_avalon_slave_0_writedata;         // mm_interconnect_0:laser_driver_avalon_slave_0_writedata -> laser_driver:avmms_writedata
	wire   [2:0] mm_interconnect_0_laser_driver_avalon_slave_0_address;           // mm_interconnect_0:laser_driver_avalon_slave_0_address -> laser_driver:avmms_address
	wire         mm_interconnect_0_laser_driver_avalon_slave_0_chipselect;        // mm_interconnect_0:laser_driver_avalon_slave_0_chipselect -> laser_driver:avmms_cs
	wire         mm_interconnect_0_laser_driver_avalon_slave_0_write;             // mm_interconnect_0:laser_driver_avalon_slave_0_write -> laser_driver:avmms_write
	wire         mm_interconnect_0_laser_driver_avalon_slave_0_read;              // mm_interconnect_0:laser_driver_avalon_slave_0_read -> laser_driver:avmms_read
	wire  [31:0] mm_interconnect_0_laser_driver_avalon_slave_0_readdata;          // laser_driver:avmms_readdata -> mm_interconnect_0:laser_driver_avalon_slave_0_readdata
	wire  [31:0] mm_interconnect_0_spi_tdc_avalon_slave_writedata;                // mm_interconnect_0:spi_tdc_avalon_slave_writedata -> spi_tdc:avmm_writedata
	wire   [1:0] mm_interconnect_0_spi_tdc_avalon_slave_address;                  // mm_interconnect_0:spi_tdc_avalon_slave_address -> spi_tdc:avmm_addr
	wire         mm_interconnect_0_spi_tdc_avalon_slave_chipselect;               // mm_interconnect_0:spi_tdc_avalon_slave_chipselect -> spi_tdc:avmm_cs
	wire         mm_interconnect_0_spi_tdc_avalon_slave_write;                    // mm_interconnect_0:spi_tdc_avalon_slave_write -> spi_tdc:avmm_write
	wire         mm_interconnect_0_spi_tdc_avalon_slave_read;                     // mm_interconnect_0:spi_tdc_avalon_slave_read -> spi_tdc:avmm_read
	wire  [31:0] mm_interconnect_0_spi_tdc_avalon_slave_readdata;                 // spi_tdc:avmm_readdata -> mm_interconnect_0:spi_tdc_avalon_slave_readdata
	wire  [31:0] mm_interconnect_0_pulse_generator_avalon_slave_writedata;        // mm_interconnect_0:pulse_generator_avalon_slave_writedata -> pulse_generator:avmm_writedata
	wire   [2:0] mm_interconnect_0_pulse_generator_avalon_slave_address;          // mm_interconnect_0:pulse_generator_avalon_slave_address -> pulse_generator:avmm_addr
	wire         mm_interconnect_0_pulse_generator_avalon_slave_chipselect;       // mm_interconnect_0:pulse_generator_avalon_slave_chipselect -> pulse_generator:avmm_cs
	wire         mm_interconnect_0_pulse_generator_avalon_slave_write;            // mm_interconnect_0:pulse_generator_avalon_slave_write -> pulse_generator:avmm_write
	wire         mm_interconnect_0_pulse_generator_avalon_slave_read;             // mm_interconnect_0:pulse_generator_avalon_slave_read -> pulse_generator:avmm_read
	wire  [31:0] mm_interconnect_0_pulse_generator_avalon_slave_readdata;         // pulse_generator:avmm_readdata -> mm_interconnect_0:pulse_generator_avalon_slave_readdata
	wire  [31:0] mm_interconnect_0_spi_vga_avalon_slave_writedata;                // mm_interconnect_0:spi_vga_avalon_slave_writedata -> spi_vga:avmm_writedata
	wire   [1:0] mm_interconnect_0_spi_vga_avalon_slave_address;                  // mm_interconnect_0:spi_vga_avalon_slave_address -> spi_vga:avmm_addr
	wire         mm_interconnect_0_spi_vga_avalon_slave_chipselect;               // mm_interconnect_0:spi_vga_avalon_slave_chipselect -> spi_vga:avmm_cs
	wire         mm_interconnect_0_spi_vga_avalon_slave_write;                    // mm_interconnect_0:spi_vga_avalon_slave_write -> spi_vga:avmm_write
	wire         mm_interconnect_0_spi_vga_avalon_slave_read;                     // mm_interconnect_0:spi_vga_avalon_slave_read -> spi_vga:avmm_read
	wire  [31:0] mm_interconnect_0_spi_vga_avalon_slave_readdata;                 // spi_vga:avmm_readdata -> mm_interconnect_0:spi_vga_avalon_slave_readdata
	wire  [31:0] mm_interconnect_0_rs485_de_s1_writedata;                         // mm_interconnect_0:rs485_de_s1_writedata -> rs485_de:writedata
	wire   [2:0] mm_interconnect_0_rs485_de_s1_address;                           // mm_interconnect_0:rs485_de_s1_address -> rs485_de:address
	wire         mm_interconnect_0_rs485_de_s1_chipselect;                        // mm_interconnect_0:rs485_de_s1_chipselect -> rs485_de:chipselect
	wire         mm_interconnect_0_rs485_de_s1_write;                             // mm_interconnect_0:rs485_de_s1_write -> rs485_de:write_n
	wire  [31:0] mm_interconnect_0_rs485_de_s1_readdata;                          // rs485_de:readdata -> mm_interconnect_0:rs485_de_s1_readdata
	wire  [31:0] mm_interconnect_0_tdc_enable_s1_writedata;                       // mm_interconnect_0:tdc_enable_s1_writedata -> tdc_enable:writedata
	wire   [2:0] mm_interconnect_0_tdc_enable_s1_address;                         // mm_interconnect_0:tdc_enable_s1_address -> tdc_enable:address
	wire         mm_interconnect_0_tdc_enable_s1_chipselect;                      // mm_interconnect_0:tdc_enable_s1_chipselect -> tdc_enable:chipselect
	wire         mm_interconnect_0_tdc_enable_s1_write;                           // mm_interconnect_0:tdc_enable_s1_write -> tdc_enable:write_n
	wire  [31:0] mm_interconnect_0_tdc_enable_s1_readdata;                        // tdc_enable:readdata -> mm_interconnect_0:tdc_enable_s1_readdata
	wire  [15:0] mm_interconnect_0_service_timer_s1_writedata;                    // mm_interconnect_0:service_timer_s1_writedata -> service_timer:writedata
	wire   [2:0] mm_interconnect_0_service_timer_s1_address;                      // mm_interconnect_0:service_timer_s1_address -> service_timer:address
	wire         mm_interconnect_0_service_timer_s1_chipselect;                   // mm_interconnect_0:service_timer_s1_chipselect -> service_timer:chipselect
	wire         mm_interconnect_0_service_timer_s1_write;                        // mm_interconnect_0:service_timer_s1_write -> service_timer:write_n
	wire  [15:0] mm_interconnect_0_service_timer_s1_readdata;                     // service_timer:readdata -> mm_interconnect_0:service_timer_s1_readdata
	wire  [31:0] mm_interconnect_0_system_mode_s1_writedata;                      // mm_interconnect_0:system_mode_s1_writedata -> system_mode:writedata
	wire   [2:0] mm_interconnect_0_system_mode_s1_address;                        // mm_interconnect_0:system_mode_s1_address -> system_mode:address
	wire         mm_interconnect_0_system_mode_s1_chipselect;                     // mm_interconnect_0:system_mode_s1_chipselect -> system_mode:chipselect
	wire         mm_interconnect_0_system_mode_s1_write;                          // mm_interconnect_0:system_mode_s1_write -> system_mode:write_n
	wire  [31:0] mm_interconnect_0_system_mode_s1_readdata;                       // system_mode:readdata -> mm_interconnect_0:system_mode_s1_readdata
	wire  [31:0] mm_interconnect_0_amp_gain_s1_writedata;                         // mm_interconnect_0:amp_gain_s1_writedata -> amp_gain:writedata
	wire   [2:0] mm_interconnect_0_amp_gain_s1_address;                           // mm_interconnect_0:amp_gain_s1_address -> amp_gain:address
	wire         mm_interconnect_0_amp_gain_s1_chipselect;                        // mm_interconnect_0:amp_gain_s1_chipselect -> amp_gain:chipselect
	wire         mm_interconnect_0_amp_gain_s1_write;                             // mm_interconnect_0:amp_gain_s1_write -> amp_gain:write_n
	wire  [31:0] mm_interconnect_0_amp_gain_s1_readdata;                          // amp_gain:readdata -> mm_interconnect_0:amp_gain_s1_readdata
	wire   [1:0] mm_interconnect_0_apd_overcurrent_s1_address;                    // mm_interconnect_0:apd_overcurrent_s1_address -> apd_overcurrent:address
	wire  [31:0] mm_interconnect_0_apd_overcurrent_s1_readdata;                   // apd_overcurrent:readdata -> mm_interconnect_0:apd_overcurrent_s1_readdata
	wire  [31:0] mm_interconnect_0_spi_apd_avalon_slave_writedata;                // mm_interconnect_0:spi_apd_avalon_slave_writedata -> spi_apd:avmm_writedata
	wire   [1:0] mm_interconnect_0_spi_apd_avalon_slave_address;                  // mm_interconnect_0:spi_apd_avalon_slave_address -> spi_apd:avmm_addr
	wire         mm_interconnect_0_spi_apd_avalon_slave_chipselect;               // mm_interconnect_0:spi_apd_avalon_slave_chipselect -> spi_apd:avmm_cs
	wire         mm_interconnect_0_spi_apd_avalon_slave_write;                    // mm_interconnect_0:spi_apd_avalon_slave_write -> spi_apd:avmm_write
	wire         mm_interconnect_0_spi_apd_avalon_slave_read;                     // mm_interconnect_0:spi_apd_avalon_slave_read -> spi_apd:avmm_read
	wire  [31:0] mm_interconnect_0_spi_apd_avalon_slave_readdata;                 // spi_apd:avmm_readdata -> mm_interconnect_0:spi_apd_avalon_slave_readdata
	wire  [31:0] mm_interconnect_0_stepper_atten_avalon_slave_0_writedata;        // mm_interconnect_0:stepper_atten_avalon_slave_0_writedata -> stepper_atten:avs_writedata
	wire   [1:0] mm_interconnect_0_stepper_atten_avalon_slave_0_address;          // mm_interconnect_0:stepper_atten_avalon_slave_0_address -> stepper_atten:avs_address
	wire         mm_interconnect_0_stepper_atten_avalon_slave_0_chipselect;       // mm_interconnect_0:stepper_atten_avalon_slave_0_chipselect -> stepper_atten:avs_cs
	wire         mm_interconnect_0_stepper_atten_avalon_slave_0_write;            // mm_interconnect_0:stepper_atten_avalon_slave_0_write -> stepper_atten:avs_write
	wire         mm_interconnect_0_stepper_atten_avalon_slave_0_read;             // mm_interconnect_0:stepper_atten_avalon_slave_0_read -> stepper_atten:avs_read
	wire  [31:0] mm_interconnect_0_stepper_atten_avalon_slave_0_readdata;         // stepper_atten:avs_readdata -> mm_interconnect_0:stepper_atten_avalon_slave_0_readdata
	wire  [31:0] mm_interconnect_0_stepper_iris_avalon_slave_0_writedata;         // mm_interconnect_0:stepper_iris_avalon_slave_0_writedata -> stepper_iris:avs_writedata
	wire   [1:0] mm_interconnect_0_stepper_iris_avalon_slave_0_address;           // mm_interconnect_0:stepper_iris_avalon_slave_0_address -> stepper_iris:avs_address
	wire         mm_interconnect_0_stepper_iris_avalon_slave_0_chipselect;        // mm_interconnect_0:stepper_iris_avalon_slave_0_chipselect -> stepper_iris:avs_cs
	wire         mm_interconnect_0_stepper_iris_avalon_slave_0_write;             // mm_interconnect_0:stepper_iris_avalon_slave_0_write -> stepper_iris:avs_write
	wire         mm_interconnect_0_stepper_iris_avalon_slave_0_read;              // mm_interconnect_0:stepper_iris_avalon_slave_0_read -> stepper_iris:avs_read
	wire  [31:0] mm_interconnect_0_stepper_iris_avalon_slave_0_readdata;          // stepper_iris:avs_readdata -> mm_interconnect_0:stepper_iris_avalon_slave_0_readdata
	wire  [31:0] mm_interconnect_0_laser_charge_avalon_slave_0_writedata;         // mm_interconnect_0:laser_charge_avalon_slave_0_writedata -> laser_charge:avmms_writedata
	wire   [2:0] mm_interconnect_0_laser_charge_avalon_slave_0_address;           // mm_interconnect_0:laser_charge_avalon_slave_0_address -> laser_charge:avmms_address
	wire         mm_interconnect_0_laser_charge_avalon_slave_0_chipselect;        // mm_interconnect_0:laser_charge_avalon_slave_0_chipselect -> laser_charge:avmms_cs
	wire         mm_interconnect_0_laser_charge_avalon_slave_0_write;             // mm_interconnect_0:laser_charge_avalon_slave_0_write -> laser_charge:avmms_write
	wire         mm_interconnect_0_laser_charge_avalon_slave_0_read;              // mm_interconnect_0:laser_charge_avalon_slave_0_read -> laser_charge:avmms_read
	wire  [31:0] mm_interconnect_0_laser_charge_avalon_slave_0_readdata;          // laser_charge:avmms_readdata -> mm_interconnect_0:laser_charge_avalon_slave_0_readdata
	wire  [31:0] mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_writedata;  // mm_interconnect_0:tdc_start_pulse_gen_avalon_slave_0_writedata -> tdc_start_pulse_gen:avmms_writedata
	wire   [2:0] mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_address;    // mm_interconnect_0:tdc_start_pulse_gen_avalon_slave_0_address -> tdc_start_pulse_gen:avmms_address
	wire         mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_chipselect; // mm_interconnect_0:tdc_start_pulse_gen_avalon_slave_0_chipselect -> tdc_start_pulse_gen:avmms_cs
	wire         mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_write;      // mm_interconnect_0:tdc_start_pulse_gen_avalon_slave_0_write -> tdc_start_pulse_gen:avmms_write
	wire         mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_read;       // mm_interconnect_0:tdc_start_pulse_gen_avalon_slave_0_read -> tdc_start_pulse_gen:avmms_read
	wire  [31:0] mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_readdata;   // tdc_start_pulse_gen:avmms_readdata -> mm_interconnect_0:tdc_start_pulse_gen_avalon_slave_0_readdata
	wire  [31:0] mm_interconnect_0_sample_recorder_avalon_slave_writedata;        // mm_interconnect_0:sample_recorder_avalon_slave_writedata -> sample_recorder:avsc_writedata
	wire   [3:0] mm_interconnect_0_sample_recorder_avalon_slave_address;          // mm_interconnect_0:sample_recorder_avalon_slave_address -> sample_recorder:avsc_addr
	wire         mm_interconnect_0_sample_recorder_avalon_slave_chipselect;       // mm_interconnect_0:sample_recorder_avalon_slave_chipselect -> sample_recorder:avsc_cs
	wire         mm_interconnect_0_sample_recorder_avalon_slave_write;            // mm_interconnect_0:sample_recorder_avalon_slave_write -> sample_recorder:avsc_write
	wire         mm_interconnect_0_sample_recorder_avalon_slave_read;             // mm_interconnect_0:sample_recorder_avalon_slave_read -> sample_recorder:avsc_read
	wire  [31:0] mm_interconnect_0_sample_recorder_avalon_slave_readdata;         // sample_recorder:avsc_readdata -> mm_interconnect_0:sample_recorder_avalon_slave_readdata
	wire   [5:0] mm_interconnect_0_sample_recorder_avalon_slave_1_address;        // mm_interconnect_0:sample_recorder_avalon_slave_1_address -> sample_recorder:avsd_addr
	wire         mm_interconnect_0_sample_recorder_avalon_slave_1_chipselect;     // mm_interconnect_0:sample_recorder_avalon_slave_1_chipselect -> sample_recorder:avsd_cs
	wire         mm_interconnect_0_sample_recorder_avalon_slave_1_read;           // mm_interconnect_0:sample_recorder_avalon_slave_1_read -> sample_recorder:avsd_read
	wire  [31:0] mm_interconnect_0_sample_recorder_avalon_slave_1_readdata;       // sample_recorder:avsd_readdata -> mm_interconnect_0:sample_recorder_avalon_slave_1_readdata
	wire         irq_mapper_receiver0_irq;                                        // sys_timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                        // pc_uart:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                        // service_timer:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_d_irq_irq;                                                   // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset]
	wire         rst_controller_reset_out_reset_req;                              // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                               // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [amp_gain:reset_n, apd_overcurrent:reset_n, i2c_port:reset_n, laser_charge:avmms_reset, laser_driver:avmms_reset, leds_port:reset_n, mm_interconnect_0:ram_cpu_reset1_reset_bridge_in_reset_reset, pc_uart:reset_n, pulse_generator:avmm_reset, ram_cpu:reset, rs485_de:reset_n, rst_translator_001:in_reset, sample_recorder:mm_reset, service_timer:reset_n, spi_apd:avmm_reset, spi_tdc:avmm_reset, spi_vga:avmm_reset, stepper_atten:avs_reset, stepper_iris:avs_reset, sys_id:reset_n, sys_timer:reset_n, system_mode:reset_n, tdc_enable:reset_n, tdc_start_pulse_gen:avmms_reset]
	wire         rst_controller_001_reset_out_reset_req;                          // rst_controller_001:reset_req -> [ram_cpu:reset_req, rst_translator_001:reset_req_in]

	rangefinder_sopc_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	rangefinder_sopc_ram_cpu ram_cpu (
		.address     (mm_interconnect_0_ram_cpu_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_ram_cpu_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_ram_cpu_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_ram_cpu_s1_write),      //       .write
		.readdata    (mm_interconnect_0_ram_cpu_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_ram_cpu_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_ram_cpu_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_ram_cpu_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_ram_cpu_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_ram_cpu_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_ram_cpu_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_ram_cpu_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_ram_cpu_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_ram_cpu_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                                 //   clk1.clk
		.reset       (rst_controller_001_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req)   //       .reset_req
	);

	rangefinder_sopc_sys_id sys_id (
		.clock    (clk_clk),                                         //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),             //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	rangefinder_sopc_sys_timer sys_timer (
		.clk           (clk_clk),                                   //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),       //         reset.reset_n
		.address       (mm_interconnect_0_sys_timer_s1_address),    //            s1.address
		.writedata     (mm_interconnect_0_sys_timer_s1_writedata),  //              .writedata
		.readdata      (mm_interconnect_0_sys_timer_s1_readdata),   //              .readdata
		.chipselect    (mm_interconnect_0_sys_timer_s1_chipselect), //              .chipselect
		.write_n       (~mm_interconnect_0_sys_timer_s1_write),     //              .write_n
		.irq           (irq_mapper_receiver0_irq),                  //           irq.irq
		.timeout_pulse (sys_timer_export)                           // external_port.export
	);

	rangefinder_sopc_pc_uart pc_uart (
		.clk           (clk_clk),                                    //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address       (mm_interconnect_0_pc_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_pc_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_pc_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_pc_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_pc_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_pc_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_pc_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                           //                    .dataavailable
		.readyfordata  (),                                           //                    .readyfordata
		.rxd           (pc_uart_rxd),                                // external_connection.export
		.txd           (pc_uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver1_irq)                    //                 irq.irq
	);

	rangefinder_sopc_leds_port leds_port (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_leds_port_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_port_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_port_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_port_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_port_s1_readdata),   //                    .readdata
		.out_port   (leds_port_export)                           // external_connection.export
	);

	rangefinder_sopc_i2c_port i2c_port (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_i2c_port_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_i2c_port_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_i2c_port_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_i2c_port_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_i2c_port_s1_readdata),   //                    .readdata
		.bidir_port (i2c_port_export)                           // external_connection.export
	);

	laser_driver laser_driver (
		.avmms_cs        (mm_interconnect_0_laser_driver_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avmms_address   (mm_interconnect_0_laser_driver_avalon_slave_0_address),    //               .address
		.avmms_write     (mm_interconnect_0_laser_driver_avalon_slave_0_write),      //               .write
		.avmms_writedata (mm_interconnect_0_laser_driver_avalon_slave_0_writedata),  //               .writedata
		.avmms_read      (mm_interconnect_0_laser_driver_avalon_slave_0_read),       //               .read
		.avmms_readdata  (mm_interconnect_0_laser_driver_avalon_slave_0_readdata),   //               .readdata
		.ref_clk         (laser_driver_ref_clk),                                     //    conduit_end.ref_clk
		.driver_mod_en   (laser_driver_driver_enable),                               //               .driver_enable
		.laser_en        (laser_driver_laser),                                       //               .laser
		.comparator      (laser_driver_comparator),                                  //               .comparator
		.avmms_clk       (clk_clk),                                                  //     clock_sink.clk
		.avmms_reset     (rst_controller_001_reset_out_reset)                        //     reset_sink.reset
	);

	spi_controller spi_tdc (
		.avmm_reset     (rst_controller_001_reset_out_reset),                //   reset_sink.reset
		.avmm_clk       (clk_clk),                                           //   clock_sink.clk
		.spi_clk        (spi_tdc_master_clk),                                //  conduit_end.master_clk
		.spi_cs_n       (spi_tdc_master_csn),                                //             .master_csn
		.spi_mosi       (spi_tdc_master_mosi),                               //             .master_mosi
		.spi_miso       (spi_tdc_master_miso),                               //             .master_miso
		.avmm_addr      (mm_interconnect_0_spi_tdc_avalon_slave_address),    // avalon_slave.address
		.avmm_cs        (mm_interconnect_0_spi_tdc_avalon_slave_chipselect), //             .chipselect
		.avmm_write     (mm_interconnect_0_spi_tdc_avalon_slave_write),      //             .write
		.avmm_writedata (mm_interconnect_0_spi_tdc_avalon_slave_writedata),  //             .writedata
		.avmm_read      (mm_interconnect_0_spi_tdc_avalon_slave_read),       //             .read
		.avmm_readdata  (mm_interconnect_0_spi_tdc_avalon_slave_readdata)    //             .readdata
	);

	test_pulse_generator pulse_generator (
		.avmm_reset     (rst_controller_001_reset_out_reset),                        //   reset_sink.reset
		.avmm_clk       (clk_clk),                                                   //   clock_sink.clk
		.start_pulse    (pulse_generator_start_pulse),                               //  conduit_end.start_pulse
		.stop_pulse     (pulse_generator_stop_pulse),                                //             .stop_pulse
		.avmm_cs        (mm_interconnect_0_pulse_generator_avalon_slave_chipselect), // avalon_slave.chipselect
		.avmm_addr      (mm_interconnect_0_pulse_generator_avalon_slave_address),    //             .address
		.avmm_write     (mm_interconnect_0_pulse_generator_avalon_slave_write),      //             .write
		.avmm_writedata (mm_interconnect_0_pulse_generator_avalon_slave_writedata),  //             .writedata
		.avmm_read      (mm_interconnect_0_pulse_generator_avalon_slave_read),       //             .read
		.avmm_readdata  (mm_interconnect_0_pulse_generator_avalon_slave_readdata)    //             .readdata
	);

	spi_controller spi_vga (
		.avmm_reset     (rst_controller_001_reset_out_reset),                //   reset_sink.reset
		.avmm_clk       (clk_clk),                                           //   clock_sink.clk
		.spi_clk        (spi_vga_master_clk),                                //  conduit_end.master_clk
		.spi_cs_n       (spi_vga_master_csn),                                //             .master_csn
		.spi_mosi       (spi_vga_master_mosi),                               //             .master_mosi
		.spi_miso       (spi_vga_master_miso),                               //             .master_miso
		.avmm_addr      (mm_interconnect_0_spi_vga_avalon_slave_address),    // avalon_slave.address
		.avmm_cs        (mm_interconnect_0_spi_vga_avalon_slave_chipselect), //             .chipselect
		.avmm_write     (mm_interconnect_0_spi_vga_avalon_slave_write),      //             .write
		.avmm_writedata (mm_interconnect_0_spi_vga_avalon_slave_writedata),  //             .writedata
		.avmm_read      (mm_interconnect_0_spi_vga_avalon_slave_read),       //             .read
		.avmm_readdata  (mm_interconnect_0_spi_vga_avalon_slave_readdata)    //             .readdata
	);

	rangefinder_sopc_rs485_de rs485_de (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_rs485_de_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_rs485_de_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_rs485_de_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_rs485_de_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_rs485_de_s1_readdata),   //                    .readdata
		.out_port   (rs485_de_export)                           // external_connection.export
	);

	rangefinder_sopc_rs485_de tdc_enable (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_tdc_enable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tdc_enable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tdc_enable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tdc_enable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tdc_enable_s1_readdata),   //                    .readdata
		.out_port   (tdc_enable_export)                           // external_connection.export
	);

	rangefinder_sopc_service_timer service_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_service_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_service_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_service_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_service_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_service_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                       //   irq.irq
	);

	spi_controller spi_apd (
		.avmm_reset     (rst_controller_001_reset_out_reset),                //   reset_sink.reset
		.avmm_clk       (clk_clk),                                           //   clock_sink.clk
		.spi_clk        (spi_apd_master_clk),                                //  conduit_end.master_clk
		.spi_cs_n       (spi_apd_master_csn),                                //             .master_csn
		.spi_mosi       (spi_apd_master_mosi),                               //             .master_mosi
		.spi_miso       (spi_apd_master_miso),                               //             .master_miso
		.avmm_addr      (mm_interconnect_0_spi_apd_avalon_slave_address),    // avalon_slave.address
		.avmm_cs        (mm_interconnect_0_spi_apd_avalon_slave_chipselect), //             .chipselect
		.avmm_write     (mm_interconnect_0_spi_apd_avalon_slave_write),      //             .write
		.avmm_writedata (mm_interconnect_0_spi_apd_avalon_slave_writedata),  //             .writedata
		.avmm_read      (mm_interconnect_0_spi_apd_avalon_slave_read),       //             .read
		.avmm_readdata  (mm_interconnect_0_spi_apd_avalon_slave_readdata)    //             .readdata
	);

	rangefinder_sopc_rs485_de system_mode (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_system_mode_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_system_mode_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_system_mode_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_system_mode_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_system_mode_s1_readdata),   //                    .readdata
		.out_port   (system_mode_export)                           // external_connection.export
	);

	rangefinder_sopc_rs485_de amp_gain (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_amp_gain_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_amp_gain_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_amp_gain_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_amp_gain_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_amp_gain_s1_readdata),   //                    .readdata
		.out_port   (amp_gain_export)                           // external_connection.export
	);

	rangefinder_sopc_apd_overcurrent apd_overcurrent (
		.clk      (clk_clk),                                       //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_apd_overcurrent_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_apd_overcurrent_s1_readdata), //                    .readdata
		.in_port  (apd_overcurrent_export)                         // external_connection.export
	);

	stepper_controller stepper_atten (
		.avs_cs        (mm_interconnect_0_stepper_atten_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avs_address   (mm_interconnect_0_stepper_atten_avalon_slave_0_address),    //               .address
		.avs_write     (mm_interconnect_0_stepper_atten_avalon_slave_0_write),      //               .write
		.avs_writedata (mm_interconnect_0_stepper_atten_avalon_slave_0_writedata),  //               .writedata
		.avs_read      (mm_interconnect_0_stepper_atten_avalon_slave_0_read),       //               .read
		.avs_readdata  (mm_interconnect_0_stepper_atten_avalon_slave_0_readdata),   //               .readdata
		.avs_clk       (clk_clk),                                                   //     clock_sink.clk
		.avs_reset     (rst_controller_001_reset_out_reset),                        //     reset_sink.reset
		.dir           (atten_motor_dir),                                           //    conduit_end.motor_dir
		.step          (atten_motor_step),                                          //               .motor_step
		.en            (atten_motor_en)                                             //               .motor_en
	);

	stepper_controller stepper_iris (
		.avs_cs        (mm_interconnect_0_stepper_iris_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avs_address   (mm_interconnect_0_stepper_iris_avalon_slave_0_address),    //               .address
		.avs_write     (mm_interconnect_0_stepper_iris_avalon_slave_0_write),      //               .write
		.avs_writedata (mm_interconnect_0_stepper_iris_avalon_slave_0_writedata),  //               .writedata
		.avs_read      (mm_interconnect_0_stepper_iris_avalon_slave_0_read),       //               .read
		.avs_readdata  (mm_interconnect_0_stepper_iris_avalon_slave_0_readdata),   //               .readdata
		.avs_clk       (clk_clk),                                                  //     clock_sink.clk
		.avs_reset     (rst_controller_001_reset_out_reset),                       //     reset_sink.reset
		.dir           (iris_motor_dir),                                           //    conduit_end.motor_dir
		.step          (iris_motor_step),                                          //               .motor_step
		.en            (iris_motor_en)                                             //               .motor_en
	);

	laser_driver laser_charge (
		.avmms_cs        (mm_interconnect_0_laser_charge_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avmms_address   (mm_interconnect_0_laser_charge_avalon_slave_0_address),    //               .address
		.avmms_write     (mm_interconnect_0_laser_charge_avalon_slave_0_write),      //               .write
		.avmms_writedata (mm_interconnect_0_laser_charge_avalon_slave_0_writedata),  //               .writedata
		.avmms_read      (mm_interconnect_0_laser_charge_avalon_slave_0_read),       //               .read
		.avmms_readdata  (mm_interconnect_0_laser_charge_avalon_slave_0_readdata),   //               .readdata
		.ref_clk         (laser_charge_ref_clk),                                     //    conduit_end.ref_clk
		.driver_mod_en   (laser_charge_driver_enable),                               //               .driver_enable
		.laser_en        (laser_charge_laser),                                       //               .laser
		.comparator      (laser_charge_comparator),                                  //               .comparator
		.avmms_clk       (clk_clk),                                                  //     clock_sink.clk
		.avmms_reset     (rst_controller_001_reset_out_reset)                        //     reset_sink.reset
	);

	laser_driver tdc_start_pulse_gen (
		.avmms_cs        (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.avmms_address   (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_address),    //               .address
		.avmms_write     (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_write),      //               .write
		.avmms_writedata (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_writedata),  //               .writedata
		.avmms_read      (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_read),       //               .read
		.avmms_readdata  (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_readdata),   //               .readdata
		.ref_clk         (tdc_start_pulse_gen_ref_clk),                                     //    conduit_end.ref_clk
		.driver_mod_en   (tdc_start_pulse_gen_driver_enable),                               //               .driver_enable
		.laser_en        (tdc_start_pulse_gen_laser),                                       //               .laser
		.comparator      (tdc_start_pulse_gen_comparator),                                  //               .comparator
		.avmms_clk       (clk_clk),                                                         //     clock_sink.clk
		.avmms_reset     (rst_controller_001_reset_out_reset)                               //     reset_sink.reset
	);

	sample_recorder sample_recorder (
		.mm_clk         (clk_clk),                                                     //     clock_sink.clk
		.mm_reset       (rst_controller_001_reset_out_reset),                          //     reset_sink.reset
		.avsc_cs        (mm_interconnect_0_sample_recorder_avalon_slave_chipselect),   //   avalon_slave.chipselect
		.avsc_addr      (mm_interconnect_0_sample_recorder_avalon_slave_address),      //               .address
		.avsc_write     (mm_interconnect_0_sample_recorder_avalon_slave_write),        //               .write
		.avsc_writedata (mm_interconnect_0_sample_recorder_avalon_slave_writedata),    //               .writedata
		.avsc_read      (mm_interconnect_0_sample_recorder_avalon_slave_read),         //               .read
		.avsc_readdata  (mm_interconnect_0_sample_recorder_avalon_slave_readdata),     //               .readdata
		.avsd_cs        (mm_interconnect_0_sample_recorder_avalon_slave_1_chipselect), // avalon_slave_1.chipselect
		.avsd_addr      (mm_interconnect_0_sample_recorder_avalon_slave_1_address),    //               .address
		.avsd_read      (mm_interconnect_0_sample_recorder_avalon_slave_1_read),       //               .read
		.avsd_readdata  (mm_interconnect_0_sample_recorder_avalon_slave_1_readdata),   //               .readdata
		.adc_clk        (adc_clk_clk),                                                 //   clock_sink_1.clk
		.adc_data       (adc_data_adc_data),                                           //    conduit_end.adc_data
		.comparator     (adc_data_comparator)                                          //               .comparator
	);

	rangefinder_sopc_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                   (clk_clk),                                                         //                              clk_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                  //    cpu_reset_n_reset_bridge_in_reset.reset
		.ram_cpu_reset1_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                              // ram_cpu_reset1_reset_bridge_in_reset.reset
		.cpu_data_master_address                       (cpu_data_master_address),                                         //                      cpu_data_master.address
		.cpu_data_master_waitrequest                   (cpu_data_master_waitrequest),                                     //                                     .waitrequest
		.cpu_data_master_byteenable                    (cpu_data_master_byteenable),                                      //                                     .byteenable
		.cpu_data_master_read                          (cpu_data_master_read),                                            //                                     .read
		.cpu_data_master_readdata                      (cpu_data_master_readdata),                                        //                                     .readdata
		.cpu_data_master_readdatavalid                 (cpu_data_master_readdatavalid),                                   //                                     .readdatavalid
		.cpu_data_master_write                         (cpu_data_master_write),                                           //                                     .write
		.cpu_data_master_writedata                     (cpu_data_master_writedata),                                       //                                     .writedata
		.cpu_data_master_debugaccess                   (cpu_data_master_debugaccess),                                     //                                     .debugaccess
		.cpu_instruction_master_address                (cpu_instruction_master_address),                                  //               cpu_instruction_master.address
		.cpu_instruction_master_waitrequest            (cpu_instruction_master_waitrequest),                              //                                     .waitrequest
		.cpu_instruction_master_read                   (cpu_instruction_master_read),                                     //                                     .read
		.cpu_instruction_master_readdata               (cpu_instruction_master_readdata),                                 //                                     .readdata
		.cpu_instruction_master_readdatavalid          (cpu_instruction_master_readdatavalid),                            //                                     .readdatavalid
		.amp_gain_s1_address                           (mm_interconnect_0_amp_gain_s1_address),                           //                          amp_gain_s1.address
		.amp_gain_s1_write                             (mm_interconnect_0_amp_gain_s1_write),                             //                                     .write
		.amp_gain_s1_readdata                          (mm_interconnect_0_amp_gain_s1_readdata),                          //                                     .readdata
		.amp_gain_s1_writedata                         (mm_interconnect_0_amp_gain_s1_writedata),                         //                                     .writedata
		.amp_gain_s1_chipselect                        (mm_interconnect_0_amp_gain_s1_chipselect),                        //                                     .chipselect
		.apd_overcurrent_s1_address                    (mm_interconnect_0_apd_overcurrent_s1_address),                    //                   apd_overcurrent_s1.address
		.apd_overcurrent_s1_readdata                   (mm_interconnect_0_apd_overcurrent_s1_readdata),                   //                                     .readdata
		.cpu_jtag_debug_module_address                 (mm_interconnect_0_cpu_jtag_debug_module_address),                 //                cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                   (mm_interconnect_0_cpu_jtag_debug_module_write),                   //                                     .write
		.cpu_jtag_debug_module_read                    (mm_interconnect_0_cpu_jtag_debug_module_read),                    //                                     .read
		.cpu_jtag_debug_module_readdata                (mm_interconnect_0_cpu_jtag_debug_module_readdata),                //                                     .readdata
		.cpu_jtag_debug_module_writedata               (mm_interconnect_0_cpu_jtag_debug_module_writedata),               //                                     .writedata
		.cpu_jtag_debug_module_byteenable              (mm_interconnect_0_cpu_jtag_debug_module_byteenable),              //                                     .byteenable
		.cpu_jtag_debug_module_waitrequest             (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),             //                                     .waitrequest
		.cpu_jtag_debug_module_debugaccess             (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),             //                                     .debugaccess
		.i2c_port_s1_address                           (mm_interconnect_0_i2c_port_s1_address),                           //                          i2c_port_s1.address
		.i2c_port_s1_write                             (mm_interconnect_0_i2c_port_s1_write),                             //                                     .write
		.i2c_port_s1_readdata                          (mm_interconnect_0_i2c_port_s1_readdata),                          //                                     .readdata
		.i2c_port_s1_writedata                         (mm_interconnect_0_i2c_port_s1_writedata),                         //                                     .writedata
		.i2c_port_s1_chipselect                        (mm_interconnect_0_i2c_port_s1_chipselect),                        //                                     .chipselect
		.laser_charge_avalon_slave_0_address           (mm_interconnect_0_laser_charge_avalon_slave_0_address),           //          laser_charge_avalon_slave_0.address
		.laser_charge_avalon_slave_0_write             (mm_interconnect_0_laser_charge_avalon_slave_0_write),             //                                     .write
		.laser_charge_avalon_slave_0_read              (mm_interconnect_0_laser_charge_avalon_slave_0_read),              //                                     .read
		.laser_charge_avalon_slave_0_readdata          (mm_interconnect_0_laser_charge_avalon_slave_0_readdata),          //                                     .readdata
		.laser_charge_avalon_slave_0_writedata         (mm_interconnect_0_laser_charge_avalon_slave_0_writedata),         //                                     .writedata
		.laser_charge_avalon_slave_0_chipselect        (mm_interconnect_0_laser_charge_avalon_slave_0_chipselect),        //                                     .chipselect
		.laser_driver_avalon_slave_0_address           (mm_interconnect_0_laser_driver_avalon_slave_0_address),           //          laser_driver_avalon_slave_0.address
		.laser_driver_avalon_slave_0_write             (mm_interconnect_0_laser_driver_avalon_slave_0_write),             //                                     .write
		.laser_driver_avalon_slave_0_read              (mm_interconnect_0_laser_driver_avalon_slave_0_read),              //                                     .read
		.laser_driver_avalon_slave_0_readdata          (mm_interconnect_0_laser_driver_avalon_slave_0_readdata),          //                                     .readdata
		.laser_driver_avalon_slave_0_writedata         (mm_interconnect_0_laser_driver_avalon_slave_0_writedata),         //                                     .writedata
		.laser_driver_avalon_slave_0_chipselect        (mm_interconnect_0_laser_driver_avalon_slave_0_chipselect),        //                                     .chipselect
		.leds_port_s1_address                          (mm_interconnect_0_leds_port_s1_address),                          //                         leds_port_s1.address
		.leds_port_s1_write                            (mm_interconnect_0_leds_port_s1_write),                            //                                     .write
		.leds_port_s1_readdata                         (mm_interconnect_0_leds_port_s1_readdata),                         //                                     .readdata
		.leds_port_s1_writedata                        (mm_interconnect_0_leds_port_s1_writedata),                        //                                     .writedata
		.leds_port_s1_chipselect                       (mm_interconnect_0_leds_port_s1_chipselect),                       //                                     .chipselect
		.pc_uart_s1_address                            (mm_interconnect_0_pc_uart_s1_address),                            //                           pc_uart_s1.address
		.pc_uart_s1_write                              (mm_interconnect_0_pc_uart_s1_write),                              //                                     .write
		.pc_uart_s1_read                               (mm_interconnect_0_pc_uart_s1_read),                               //                                     .read
		.pc_uart_s1_readdata                           (mm_interconnect_0_pc_uart_s1_readdata),                           //                                     .readdata
		.pc_uart_s1_writedata                          (mm_interconnect_0_pc_uart_s1_writedata),                          //                                     .writedata
		.pc_uart_s1_begintransfer                      (mm_interconnect_0_pc_uart_s1_begintransfer),                      //                                     .begintransfer
		.pc_uart_s1_chipselect                         (mm_interconnect_0_pc_uart_s1_chipselect),                         //                                     .chipselect
		.pulse_generator_avalon_slave_address          (mm_interconnect_0_pulse_generator_avalon_slave_address),          //         pulse_generator_avalon_slave.address
		.pulse_generator_avalon_slave_write            (mm_interconnect_0_pulse_generator_avalon_slave_write),            //                                     .write
		.pulse_generator_avalon_slave_read             (mm_interconnect_0_pulse_generator_avalon_slave_read),             //                                     .read
		.pulse_generator_avalon_slave_readdata         (mm_interconnect_0_pulse_generator_avalon_slave_readdata),         //                                     .readdata
		.pulse_generator_avalon_slave_writedata        (mm_interconnect_0_pulse_generator_avalon_slave_writedata),        //                                     .writedata
		.pulse_generator_avalon_slave_chipselect       (mm_interconnect_0_pulse_generator_avalon_slave_chipselect),       //                                     .chipselect
		.ram_cpu_s1_address                            (mm_interconnect_0_ram_cpu_s1_address),                            //                           ram_cpu_s1.address
		.ram_cpu_s1_write                              (mm_interconnect_0_ram_cpu_s1_write),                              //                                     .write
		.ram_cpu_s1_readdata                           (mm_interconnect_0_ram_cpu_s1_readdata),                           //                                     .readdata
		.ram_cpu_s1_writedata                          (mm_interconnect_0_ram_cpu_s1_writedata),                          //                                     .writedata
		.ram_cpu_s1_byteenable                         (mm_interconnect_0_ram_cpu_s1_byteenable),                         //                                     .byteenable
		.ram_cpu_s1_chipselect                         (mm_interconnect_0_ram_cpu_s1_chipselect),                         //                                     .chipselect
		.ram_cpu_s1_clken                              (mm_interconnect_0_ram_cpu_s1_clken),                              //                                     .clken
		.ram_cpu_s2_address                            (mm_interconnect_0_ram_cpu_s2_address),                            //                           ram_cpu_s2.address
		.ram_cpu_s2_write                              (mm_interconnect_0_ram_cpu_s2_write),                              //                                     .write
		.ram_cpu_s2_readdata                           (mm_interconnect_0_ram_cpu_s2_readdata),                           //                                     .readdata
		.ram_cpu_s2_writedata                          (mm_interconnect_0_ram_cpu_s2_writedata),                          //                                     .writedata
		.ram_cpu_s2_byteenable                         (mm_interconnect_0_ram_cpu_s2_byteenable),                         //                                     .byteenable
		.ram_cpu_s2_chipselect                         (mm_interconnect_0_ram_cpu_s2_chipselect),                         //                                     .chipselect
		.ram_cpu_s2_clken                              (mm_interconnect_0_ram_cpu_s2_clken),                              //                                     .clken
		.rs485_de_s1_address                           (mm_interconnect_0_rs485_de_s1_address),                           //                          rs485_de_s1.address
		.rs485_de_s1_write                             (mm_interconnect_0_rs485_de_s1_write),                             //                                     .write
		.rs485_de_s1_readdata                          (mm_interconnect_0_rs485_de_s1_readdata),                          //                                     .readdata
		.rs485_de_s1_writedata                         (mm_interconnect_0_rs485_de_s1_writedata),                         //                                     .writedata
		.rs485_de_s1_chipselect                        (mm_interconnect_0_rs485_de_s1_chipselect),                        //                                     .chipselect
		.sample_recorder_avalon_slave_address          (mm_interconnect_0_sample_recorder_avalon_slave_address),          //         sample_recorder_avalon_slave.address
		.sample_recorder_avalon_slave_write            (mm_interconnect_0_sample_recorder_avalon_slave_write),            //                                     .write
		.sample_recorder_avalon_slave_read             (mm_interconnect_0_sample_recorder_avalon_slave_read),             //                                     .read
		.sample_recorder_avalon_slave_readdata         (mm_interconnect_0_sample_recorder_avalon_slave_readdata),         //                                     .readdata
		.sample_recorder_avalon_slave_writedata        (mm_interconnect_0_sample_recorder_avalon_slave_writedata),        //                                     .writedata
		.sample_recorder_avalon_slave_chipselect       (mm_interconnect_0_sample_recorder_avalon_slave_chipselect),       //                                     .chipselect
		.sample_recorder_avalon_slave_1_address        (mm_interconnect_0_sample_recorder_avalon_slave_1_address),        //       sample_recorder_avalon_slave_1.address
		.sample_recorder_avalon_slave_1_read           (mm_interconnect_0_sample_recorder_avalon_slave_1_read),           //                                     .read
		.sample_recorder_avalon_slave_1_readdata       (mm_interconnect_0_sample_recorder_avalon_slave_1_readdata),       //                                     .readdata
		.sample_recorder_avalon_slave_1_chipselect     (mm_interconnect_0_sample_recorder_avalon_slave_1_chipselect),     //                                     .chipselect
		.service_timer_s1_address                      (mm_interconnect_0_service_timer_s1_address),                      //                     service_timer_s1.address
		.service_timer_s1_write                        (mm_interconnect_0_service_timer_s1_write),                        //                                     .write
		.service_timer_s1_readdata                     (mm_interconnect_0_service_timer_s1_readdata),                     //                                     .readdata
		.service_timer_s1_writedata                    (mm_interconnect_0_service_timer_s1_writedata),                    //                                     .writedata
		.service_timer_s1_chipselect                   (mm_interconnect_0_service_timer_s1_chipselect),                   //                                     .chipselect
		.spi_apd_avalon_slave_address                  (mm_interconnect_0_spi_apd_avalon_slave_address),                  //                 spi_apd_avalon_slave.address
		.spi_apd_avalon_slave_write                    (mm_interconnect_0_spi_apd_avalon_slave_write),                    //                                     .write
		.spi_apd_avalon_slave_read                     (mm_interconnect_0_spi_apd_avalon_slave_read),                     //                                     .read
		.spi_apd_avalon_slave_readdata                 (mm_interconnect_0_spi_apd_avalon_slave_readdata),                 //                                     .readdata
		.spi_apd_avalon_slave_writedata                (mm_interconnect_0_spi_apd_avalon_slave_writedata),                //                                     .writedata
		.spi_apd_avalon_slave_chipselect               (mm_interconnect_0_spi_apd_avalon_slave_chipselect),               //                                     .chipselect
		.spi_tdc_avalon_slave_address                  (mm_interconnect_0_spi_tdc_avalon_slave_address),                  //                 spi_tdc_avalon_slave.address
		.spi_tdc_avalon_slave_write                    (mm_interconnect_0_spi_tdc_avalon_slave_write),                    //                                     .write
		.spi_tdc_avalon_slave_read                     (mm_interconnect_0_spi_tdc_avalon_slave_read),                     //                                     .read
		.spi_tdc_avalon_slave_readdata                 (mm_interconnect_0_spi_tdc_avalon_slave_readdata),                 //                                     .readdata
		.spi_tdc_avalon_slave_writedata                (mm_interconnect_0_spi_tdc_avalon_slave_writedata),                //                                     .writedata
		.spi_tdc_avalon_slave_chipselect               (mm_interconnect_0_spi_tdc_avalon_slave_chipselect),               //                                     .chipselect
		.spi_vga_avalon_slave_address                  (mm_interconnect_0_spi_vga_avalon_slave_address),                  //                 spi_vga_avalon_slave.address
		.spi_vga_avalon_slave_write                    (mm_interconnect_0_spi_vga_avalon_slave_write),                    //                                     .write
		.spi_vga_avalon_slave_read                     (mm_interconnect_0_spi_vga_avalon_slave_read),                     //                                     .read
		.spi_vga_avalon_slave_readdata                 (mm_interconnect_0_spi_vga_avalon_slave_readdata),                 //                                     .readdata
		.spi_vga_avalon_slave_writedata                (mm_interconnect_0_spi_vga_avalon_slave_writedata),                //                                     .writedata
		.spi_vga_avalon_slave_chipselect               (mm_interconnect_0_spi_vga_avalon_slave_chipselect),               //                                     .chipselect
		.stepper_atten_avalon_slave_0_address          (mm_interconnect_0_stepper_atten_avalon_slave_0_address),          //         stepper_atten_avalon_slave_0.address
		.stepper_atten_avalon_slave_0_write            (mm_interconnect_0_stepper_atten_avalon_slave_0_write),            //                                     .write
		.stepper_atten_avalon_slave_0_read             (mm_interconnect_0_stepper_atten_avalon_slave_0_read),             //                                     .read
		.stepper_atten_avalon_slave_0_readdata         (mm_interconnect_0_stepper_atten_avalon_slave_0_readdata),         //                                     .readdata
		.stepper_atten_avalon_slave_0_writedata        (mm_interconnect_0_stepper_atten_avalon_slave_0_writedata),        //                                     .writedata
		.stepper_atten_avalon_slave_0_chipselect       (mm_interconnect_0_stepper_atten_avalon_slave_0_chipselect),       //                                     .chipselect
		.stepper_iris_avalon_slave_0_address           (mm_interconnect_0_stepper_iris_avalon_slave_0_address),           //          stepper_iris_avalon_slave_0.address
		.stepper_iris_avalon_slave_0_write             (mm_interconnect_0_stepper_iris_avalon_slave_0_write),             //                                     .write
		.stepper_iris_avalon_slave_0_read              (mm_interconnect_0_stepper_iris_avalon_slave_0_read),              //                                     .read
		.stepper_iris_avalon_slave_0_readdata          (mm_interconnect_0_stepper_iris_avalon_slave_0_readdata),          //                                     .readdata
		.stepper_iris_avalon_slave_0_writedata         (mm_interconnect_0_stepper_iris_avalon_slave_0_writedata),         //                                     .writedata
		.stepper_iris_avalon_slave_0_chipselect        (mm_interconnect_0_stepper_iris_avalon_slave_0_chipselect),        //                                     .chipselect
		.sys_id_control_slave_address                  (mm_interconnect_0_sys_id_control_slave_address),                  //                 sys_id_control_slave.address
		.sys_id_control_slave_readdata                 (mm_interconnect_0_sys_id_control_slave_readdata),                 //                                     .readdata
		.sys_timer_s1_address                          (mm_interconnect_0_sys_timer_s1_address),                          //                         sys_timer_s1.address
		.sys_timer_s1_write                            (mm_interconnect_0_sys_timer_s1_write),                            //                                     .write
		.sys_timer_s1_readdata                         (mm_interconnect_0_sys_timer_s1_readdata),                         //                                     .readdata
		.sys_timer_s1_writedata                        (mm_interconnect_0_sys_timer_s1_writedata),                        //                                     .writedata
		.sys_timer_s1_chipselect                       (mm_interconnect_0_sys_timer_s1_chipselect),                       //                                     .chipselect
		.system_mode_s1_address                        (mm_interconnect_0_system_mode_s1_address),                        //                       system_mode_s1.address
		.system_mode_s1_write                          (mm_interconnect_0_system_mode_s1_write),                          //                                     .write
		.system_mode_s1_readdata                       (mm_interconnect_0_system_mode_s1_readdata),                       //                                     .readdata
		.system_mode_s1_writedata                      (mm_interconnect_0_system_mode_s1_writedata),                      //                                     .writedata
		.system_mode_s1_chipselect                     (mm_interconnect_0_system_mode_s1_chipselect),                     //                                     .chipselect
		.tdc_enable_s1_address                         (mm_interconnect_0_tdc_enable_s1_address),                         //                        tdc_enable_s1.address
		.tdc_enable_s1_write                           (mm_interconnect_0_tdc_enable_s1_write),                           //                                     .write
		.tdc_enable_s1_readdata                        (mm_interconnect_0_tdc_enable_s1_readdata),                        //                                     .readdata
		.tdc_enable_s1_writedata                       (mm_interconnect_0_tdc_enable_s1_writedata),                       //                                     .writedata
		.tdc_enable_s1_chipselect                      (mm_interconnect_0_tdc_enable_s1_chipselect),                      //                                     .chipselect
		.tdc_start_pulse_gen_avalon_slave_0_address    (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_address),    //   tdc_start_pulse_gen_avalon_slave_0.address
		.tdc_start_pulse_gen_avalon_slave_0_write      (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_write),      //                                     .write
		.tdc_start_pulse_gen_avalon_slave_0_read       (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_read),       //                                     .read
		.tdc_start_pulse_gen_avalon_slave_0_readdata   (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_readdata),   //                                     .readdata
		.tdc_start_pulse_gen_avalon_slave_0_writedata  (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_writedata),  //                                     .writedata
		.tdc_start_pulse_gen_avalon_slave_0_chipselect (mm_interconnect_0_tdc_start_pulse_gen_avalon_slave_0_chipselect)  //                                     .chipselect
	);

	rangefinder_sopc_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
